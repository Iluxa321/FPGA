
module debug (
	source,
	probe);	

	output	[7:0]	source;
	input	[9:0]	probe;
endmodule
