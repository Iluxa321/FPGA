// Размер в byte
`define UFM_OFFSET  32'h0
`define UFM_SIZE    32'h400
`define RAM_OFFSET  32'h20000
`define RAM_SIZE    32'h400



`define PERIPH_BASE  32'h40000
`define PERIPH_SIZE    32'h400

`define SEG_SIZE    32'h2
`define SEG         (`PERIPH_BASE + 4)

