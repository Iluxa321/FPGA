// Размер в byte
`define UFM_OFFSET  32'h0
`define UFM_SIZE    32'h400
`define RAM_OFFSET  32'h20000
`define RAM_SIZE    32'h400



